`ifndef PARAMETERS_VH
`define PARAMETERS_VH

`define PE_ROW 2
`define PE_COL 2

`define MM_HGT 2
`define MM_WDT 2

`define IM_HGT 2
`define IM_WDT 2
`define WM_HGT 2
`define WM_WDT 2
`define OM_HGT 2
`define OM_WDT 2

`endif